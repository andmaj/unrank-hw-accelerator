module unrank32 (
    input clk,
    input [31:0] num,
    input [5:0] col,
    output reg [5:0] row
);

wire [31:0] binom_table [1:32][1:32];
wire [1:32] bits [1:32];
wire [1:32] colbits;
wire [1:32] xorbits;
wire [5:0] irow;

assign colbits = bits[col];

always @ (posedge clk)
begin
    row <= irow;
end

// For 6-input LUT (Xilinx 7)

wire bit0_0;
wire bit0_1;
wire bit0;

assign bit0_0 = xorbits[1] | xorbits[3] | xorbits[5] | xorbits[7] | xorbits[9] | xorbits[11];
assign bit0_1 = xorbits[13] | xorbits[15] | xorbits[17] | xorbits[19] | xorbits[21] | xorbits[23];
assign bit0 = bit0_0 | bit0_1 | xorbits[25] | xorbits[27] | xorbits[29] | xorbits[31];

wire bit1_0;
wire bit1_1;
wire bit1;

assign bit1_0 = xorbits[2] | xorbits[3] | xorbits[6] | xorbits[7] | xorbits[10] | xorbits[11];
assign bit1_1 = xorbits[14] | xorbits[15] | xorbits[18] | xorbits[19] | xorbits[22] | xorbits[23];
assign bit1 = bit1_0 | bit1_1 | xorbits[26] | xorbits[27] | xorbits[30] | xorbits[31];

wire bit2_0;
wire bit2_1;
wire bit2;

assign bit2_0 = xorbits[4] | xorbits[5] | xorbits[6] | xorbits[7] | xorbits[12] | xorbits[13];
assign bit2_1 = xorbits[14] | xorbits[15] | xorbits[20] | xorbits[21] | xorbits[22] | xorbits[23];
assign bit2 = bit2_0 | bit2_1 | xorbits[28] | xorbits[29] | xorbits[30] | xorbits[31];

wire bit3_0;
wire bit3_1;
wire bit3;

assign bit3_0 = xorbits[8] | xorbits[9] | xorbits[10] | xorbits[11] | xorbits[12] | xorbits[13];
assign bit3_1 = xorbits[14] | xorbits[15] | xorbits[24] | xorbits[25] | xorbits[26] | xorbits[27];
assign bit3 = bit3_0 | bit3_1 | xorbits[28] | xorbits[29] | xorbits[30] | xorbits[31];

wire bit4_0;
wire bit4_1;
wire bit4;

assign bit4_0 = xorbits[16] | xorbits[17] | xorbits[18] | xorbits[19] | xorbits[20] | xorbits[21];
assign bit4_1 = xorbits[22] | xorbits[23] | xorbits[24] | xorbits[25] | xorbits[26] | xorbits[27];
assign bit4 = bit4_0 | bit4_1 | xorbits[28] | xorbits[29] | xorbits[30] | xorbits[31];

assign irow[0] = bit0;
assign irow[1] = bit1;
assign irow[2] = bit2;
assign irow[3] = bit3;
assign irow[4] = bit4;
assign irow[5] = xorbits[32];

assign xorbits[1] = 1^colbits[1];

/*
MAXBITS = 32

def factorial(n, stop=0):
	o = 1
	while n > stop:
		o *= n
		n -= 1
	return o

def choose(n, k):
	if n < k:
		return 0
	return factorial(n, stop=k) / factorial(n - k)

for col in range(1,MAXBITS+1):
	for row in range(1,MAXBITS+1):
		print('assign binom_table[%d][%d] = %d;' % (col, row, choose(row,col)))
	print('')

for col in range(1,MAXBITS+1):
	for row in range(1,MAXBITS+1):
		print('assign bits[%d][%d] = num > binom_table[%d][%d];' % (col, row, col, row))
	print('')

for row in range(2,MAXBITS+1):
	print('assign xorbits[%d] = colbits[%d]^colbits[%d];' % (row, row-1, row))

*/

// generated
assign binom_table[1][1] = 1;
assign binom_table[1][2] = 2;
assign binom_table[1][3] = 3;
assign binom_table[1][4] = 4;
assign binom_table[1][5] = 5;
assign binom_table[1][6] = 6;
assign binom_table[1][7] = 7;
assign binom_table[1][8] = 8;
assign binom_table[1][9] = 9;
assign binom_table[1][10] = 10;
assign binom_table[1][11] = 11;
assign binom_table[1][12] = 12;
assign binom_table[1][13] = 13;
assign binom_table[1][14] = 14;
assign binom_table[1][15] = 15;
assign binom_table[1][16] = 16;
assign binom_table[1][17] = 17;
assign binom_table[1][18] = 18;
assign binom_table[1][19] = 19;
assign binom_table[1][20] = 20;
assign binom_table[1][21] = 21;
assign binom_table[1][22] = 22;
assign binom_table[1][23] = 23;
assign binom_table[1][24] = 24;
assign binom_table[1][25] = 25;
assign binom_table[1][26] = 26;
assign binom_table[1][27] = 27;
assign binom_table[1][28] = 28;
assign binom_table[1][29] = 29;
assign binom_table[1][30] = 30;
assign binom_table[1][31] = 31;
assign binom_table[1][32] = 32;

assign binom_table[2][1] = 0;
assign binom_table[2][2] = 1;
assign binom_table[2][3] = 3;
assign binom_table[2][4] = 6;
assign binom_table[2][5] = 10;
assign binom_table[2][6] = 15;
assign binom_table[2][7] = 21;
assign binom_table[2][8] = 28;
assign binom_table[2][9] = 36;
assign binom_table[2][10] = 45;
assign binom_table[2][11] = 55;
assign binom_table[2][12] = 66;
assign binom_table[2][13] = 78;
assign binom_table[2][14] = 91;
assign binom_table[2][15] = 105;
assign binom_table[2][16] = 120;
assign binom_table[2][17] = 136;
assign binom_table[2][18] = 153;
assign binom_table[2][19] = 171;
assign binom_table[2][20] = 190;
assign binom_table[2][21] = 210;
assign binom_table[2][22] = 231;
assign binom_table[2][23] = 253;
assign binom_table[2][24] = 276;
assign binom_table[2][25] = 300;
assign binom_table[2][26] = 325;
assign binom_table[2][27] = 351;
assign binom_table[2][28] = 378;
assign binom_table[2][29] = 406;
assign binom_table[2][30] = 435;
assign binom_table[2][31] = 465;
assign binom_table[2][32] = 496;

assign binom_table[3][1] = 0;
assign binom_table[3][2] = 0;
assign binom_table[3][3] = 1;
assign binom_table[3][4] = 4;
assign binom_table[3][5] = 10;
assign binom_table[3][6] = 20;
assign binom_table[3][7] = 35;
assign binom_table[3][8] = 56;
assign binom_table[3][9] = 84;
assign binom_table[3][10] = 120;
assign binom_table[3][11] = 165;
assign binom_table[3][12] = 220;
assign binom_table[3][13] = 286;
assign binom_table[3][14] = 364;
assign binom_table[3][15] = 455;
assign binom_table[3][16] = 560;
assign binom_table[3][17] = 680;
assign binom_table[3][18] = 816;
assign binom_table[3][19] = 969;
assign binom_table[3][20] = 1140;
assign binom_table[3][21] = 1330;
assign binom_table[3][22] = 1540;
assign binom_table[3][23] = 1771;
assign binom_table[3][24] = 2024;
assign binom_table[3][25] = 2300;
assign binom_table[3][26] = 2600;
assign binom_table[3][27] = 2925;
assign binom_table[3][28] = 3276;
assign binom_table[3][29] = 3654;
assign binom_table[3][30] = 4060;
assign binom_table[3][31] = 4495;
assign binom_table[3][32] = 4960;

assign binom_table[4][1] = 0;
assign binom_table[4][2] = 0;
assign binom_table[4][3] = 0;
assign binom_table[4][4] = 1;
assign binom_table[4][5] = 5;
assign binom_table[4][6] = 15;
assign binom_table[4][7] = 35;
assign binom_table[4][8] = 70;
assign binom_table[4][9] = 126;
assign binom_table[4][10] = 210;
assign binom_table[4][11] = 330;
assign binom_table[4][12] = 495;
assign binom_table[4][13] = 715;
assign binom_table[4][14] = 1001;
assign binom_table[4][15] = 1365;
assign binom_table[4][16] = 1820;
assign binom_table[4][17] = 2380;
assign binom_table[4][18] = 3060;
assign binom_table[4][19] = 3876;
assign binom_table[4][20] = 4845;
assign binom_table[4][21] = 5985;
assign binom_table[4][22] = 7315;
assign binom_table[4][23] = 8855;
assign binom_table[4][24] = 10626;
assign binom_table[4][25] = 12650;
assign binom_table[4][26] = 14950;
assign binom_table[4][27] = 17550;
assign binom_table[4][28] = 20475;
assign binom_table[4][29] = 23751;
assign binom_table[4][30] = 27405;
assign binom_table[4][31] = 31465;
assign binom_table[4][32] = 35960;

assign binom_table[5][1] = 0;
assign binom_table[5][2] = 0;
assign binom_table[5][3] = 0;
assign binom_table[5][4] = 0;
assign binom_table[5][5] = 1;
assign binom_table[5][6] = 6;
assign binom_table[5][7] = 21;
assign binom_table[5][8] = 56;
assign binom_table[5][9] = 126;
assign binom_table[5][10] = 252;
assign binom_table[5][11] = 462;
assign binom_table[5][12] = 792;
assign binom_table[5][13] = 1287;
assign binom_table[5][14] = 2002;
assign binom_table[5][15] = 3003;
assign binom_table[5][16] = 4368;
assign binom_table[5][17] = 6188;
assign binom_table[5][18] = 8568;
assign binom_table[5][19] = 11628;
assign binom_table[5][20] = 15504;
assign binom_table[5][21] = 20349;
assign binom_table[5][22] = 26334;
assign binom_table[5][23] = 33649;
assign binom_table[5][24] = 42504;
assign binom_table[5][25] = 53130;
assign binom_table[5][26] = 65780;
assign binom_table[5][27] = 80730;
assign binom_table[5][28] = 98280;
assign binom_table[5][29] = 118755;
assign binom_table[5][30] = 142506;
assign binom_table[5][31] = 169911;
assign binom_table[5][32] = 201376;

assign binom_table[6][1] = 0;
assign binom_table[6][2] = 0;
assign binom_table[6][3] = 0;
assign binom_table[6][4] = 0;
assign binom_table[6][5] = 0;
assign binom_table[6][6] = 1;
assign binom_table[6][7] = 7;
assign binom_table[6][8] = 28;
assign binom_table[6][9] = 84;
assign binom_table[6][10] = 210;
assign binom_table[6][11] = 462;
assign binom_table[6][12] = 924;
assign binom_table[6][13] = 1716;
assign binom_table[6][14] = 3003;
assign binom_table[6][15] = 5005;
assign binom_table[6][16] = 8008;
assign binom_table[6][17] = 12376;
assign binom_table[6][18] = 18564;
assign binom_table[6][19] = 27132;
assign binom_table[6][20] = 38760;
assign binom_table[6][21] = 54264;
assign binom_table[6][22] = 74613;
assign binom_table[6][23] = 100947;
assign binom_table[6][24] = 134596;
assign binom_table[6][25] = 177100;
assign binom_table[6][26] = 230230;
assign binom_table[6][27] = 296010;
assign binom_table[6][28] = 376740;
assign binom_table[6][29] = 475020;
assign binom_table[6][30] = 593775;
assign binom_table[6][31] = 736281;
assign binom_table[6][32] = 906192;

assign binom_table[7][1] = 0;
assign binom_table[7][2] = 0;
assign binom_table[7][3] = 0;
assign binom_table[7][4] = 0;
assign binom_table[7][5] = 0;
assign binom_table[7][6] = 0;
assign binom_table[7][7] = 1;
assign binom_table[7][8] = 8;
assign binom_table[7][9] = 36;
assign binom_table[7][10] = 120;
assign binom_table[7][11] = 330;
assign binom_table[7][12] = 792;
assign binom_table[7][13] = 1716;
assign binom_table[7][14] = 3432;
assign binom_table[7][15] = 6435;
assign binom_table[7][16] = 11440;
assign binom_table[7][17] = 19448;
assign binom_table[7][18] = 31824;
assign binom_table[7][19] = 50388;
assign binom_table[7][20] = 77520;
assign binom_table[7][21] = 116280;
assign binom_table[7][22] = 170544;
assign binom_table[7][23] = 245157;
assign binom_table[7][24] = 346104;
assign binom_table[7][25] = 480700;
assign binom_table[7][26] = 657800;
assign binom_table[7][27] = 888030;
assign binom_table[7][28] = 1184040;
assign binom_table[7][29] = 1560780;
assign binom_table[7][30] = 2035800;
assign binom_table[7][31] = 2629575;
assign binom_table[7][32] = 3365856;

assign binom_table[8][1] = 0;
assign binom_table[8][2] = 0;
assign binom_table[8][3] = 0;
assign binom_table[8][4] = 0;
assign binom_table[8][5] = 0;
assign binom_table[8][6] = 0;
assign binom_table[8][7] = 0;
assign binom_table[8][8] = 1;
assign binom_table[8][9] = 9;
assign binom_table[8][10] = 45;
assign binom_table[8][11] = 165;
assign binom_table[8][12] = 495;
assign binom_table[8][13] = 1287;
assign binom_table[8][14] = 3003;
assign binom_table[8][15] = 6435;
assign binom_table[8][16] = 12870;
assign binom_table[8][17] = 24310;
assign binom_table[8][18] = 43758;
assign binom_table[8][19] = 75582;
assign binom_table[8][20] = 125970;
assign binom_table[8][21] = 203490;
assign binom_table[8][22] = 319770;
assign binom_table[8][23] = 490314;
assign binom_table[8][24] = 735471;
assign binom_table[8][25] = 1081575;
assign binom_table[8][26] = 1562275;
assign binom_table[8][27] = 2220075;
assign binom_table[8][28] = 3108105;
assign binom_table[8][29] = 4292145;
assign binom_table[8][30] = 5852925;
assign binom_table[8][31] = 7888725;
assign binom_table[8][32] = 10518300;

assign binom_table[9][1] = 0;
assign binom_table[9][2] = 0;
assign binom_table[9][3] = 0;
assign binom_table[9][4] = 0;
assign binom_table[9][5] = 0;
assign binom_table[9][6] = 0;
assign binom_table[9][7] = 0;
assign binom_table[9][8] = 0;
assign binom_table[9][9] = 1;
assign binom_table[9][10] = 10;
assign binom_table[9][11] = 55;
assign binom_table[9][12] = 220;
assign binom_table[9][13] = 715;
assign binom_table[9][14] = 2002;
assign binom_table[9][15] = 5005;
assign binom_table[9][16] = 11440;
assign binom_table[9][17] = 24310;
assign binom_table[9][18] = 48620;
assign binom_table[9][19] = 92378;
assign binom_table[9][20] = 167960;
assign binom_table[9][21] = 293930;
assign binom_table[9][22] = 497420;
assign binom_table[9][23] = 817190;
assign binom_table[9][24] = 1307504;
assign binom_table[9][25] = 2042975;
assign binom_table[9][26] = 3124550;
assign binom_table[9][27] = 4686825;
assign binom_table[9][28] = 6906900;
assign binom_table[9][29] = 10015005;
assign binom_table[9][30] = 14307150;
assign binom_table[9][31] = 20160075;
assign binom_table[9][32] = 28048800;

assign binom_table[10][1] = 0;
assign binom_table[10][2] = 0;
assign binom_table[10][3] = 0;
assign binom_table[10][4] = 0;
assign binom_table[10][5] = 0;
assign binom_table[10][6] = 0;
assign binom_table[10][7] = 0;
assign binom_table[10][8] = 0;
assign binom_table[10][9] = 0;
assign binom_table[10][10] = 1;
assign binom_table[10][11] = 11;
assign binom_table[10][12] = 66;
assign binom_table[10][13] = 286;
assign binom_table[10][14] = 1001;
assign binom_table[10][15] = 3003;
assign binom_table[10][16] = 8008;
assign binom_table[10][17] = 19448;
assign binom_table[10][18] = 43758;
assign binom_table[10][19] = 92378;
assign binom_table[10][20] = 184756;
assign binom_table[10][21] = 352716;
assign binom_table[10][22] = 646646;
assign binom_table[10][23] = 1144066;
assign binom_table[10][24] = 1961256;
assign binom_table[10][25] = 3268760;
assign binom_table[10][26] = 5311735;
assign binom_table[10][27] = 8436285;
assign binom_table[10][28] = 13123110;
assign binom_table[10][29] = 20030010;
assign binom_table[10][30] = 30045015;
assign binom_table[10][31] = 44352165;
assign binom_table[10][32] = 64512240;

assign binom_table[11][1] = 0;
assign binom_table[11][2] = 0;
assign binom_table[11][3] = 0;
assign binom_table[11][4] = 0;
assign binom_table[11][5] = 0;
assign binom_table[11][6] = 0;
assign binom_table[11][7] = 0;
assign binom_table[11][8] = 0;
assign binom_table[11][9] = 0;
assign binom_table[11][10] = 0;
assign binom_table[11][11] = 1;
assign binom_table[11][12] = 12;
assign binom_table[11][13] = 78;
assign binom_table[11][14] = 364;
assign binom_table[11][15] = 1365;
assign binom_table[11][16] = 4368;
assign binom_table[11][17] = 12376;
assign binom_table[11][18] = 31824;
assign binom_table[11][19] = 75582;
assign binom_table[11][20] = 167960;
assign binom_table[11][21] = 352716;
assign binom_table[11][22] = 705432;
assign binom_table[11][23] = 1352078;
assign binom_table[11][24] = 2496144;
assign binom_table[11][25] = 4457400;
assign binom_table[11][26] = 7726160;
assign binom_table[11][27] = 13037895;
assign binom_table[11][28] = 21474180;
assign binom_table[11][29] = 34597290;
assign binom_table[11][30] = 54627300;
assign binom_table[11][31] = 84672315;
assign binom_table[11][32] = 129024480;

assign binom_table[12][1] = 0;
assign binom_table[12][2] = 0;
assign binom_table[12][3] = 0;
assign binom_table[12][4] = 0;
assign binom_table[12][5] = 0;
assign binom_table[12][6] = 0;
assign binom_table[12][7] = 0;
assign binom_table[12][8] = 0;
assign binom_table[12][9] = 0;
assign binom_table[12][10] = 0;
assign binom_table[12][11] = 0;
assign binom_table[12][12] = 1;
assign binom_table[12][13] = 13;
assign binom_table[12][14] = 91;
assign binom_table[12][15] = 455;
assign binom_table[12][16] = 1820;
assign binom_table[12][17] = 6188;
assign binom_table[12][18] = 18564;
assign binom_table[12][19] = 50388;
assign binom_table[12][20] = 125970;
assign binom_table[12][21] = 293930;
assign binom_table[12][22] = 646646;
assign binom_table[12][23] = 1352078;
assign binom_table[12][24] = 2704156;
assign binom_table[12][25] = 5200300;
assign binom_table[12][26] = 9657700;
assign binom_table[12][27] = 17383860;
assign binom_table[12][28] = 30421755;
assign binom_table[12][29] = 51895935;
assign binom_table[12][30] = 86493225;
assign binom_table[12][31] = 141120525;
assign binom_table[12][32] = 225792840;

assign binom_table[13][1] = 0;
assign binom_table[13][2] = 0;
assign binom_table[13][3] = 0;
assign binom_table[13][4] = 0;
assign binom_table[13][5] = 0;
assign binom_table[13][6] = 0;
assign binom_table[13][7] = 0;
assign binom_table[13][8] = 0;
assign binom_table[13][9] = 0;
assign binom_table[13][10] = 0;
assign binom_table[13][11] = 0;
assign binom_table[13][12] = 0;
assign binom_table[13][13] = 1;
assign binom_table[13][14] = 14;
assign binom_table[13][15] = 105;
assign binom_table[13][16] = 560;
assign binom_table[13][17] = 2380;
assign binom_table[13][18] = 8568;
assign binom_table[13][19] = 27132;
assign binom_table[13][20] = 77520;
assign binom_table[13][21] = 203490;
assign binom_table[13][22] = 497420;
assign binom_table[13][23] = 1144066;
assign binom_table[13][24] = 2496144;
assign binom_table[13][25] = 5200300;
assign binom_table[13][26] = 10400600;
assign binom_table[13][27] = 20058300;
assign binom_table[13][28] = 37442160;
assign binom_table[13][29] = 67863915;
assign binom_table[13][30] = 119759850;
assign binom_table[13][31] = 206253075;
assign binom_table[13][32] = 347373600;

assign binom_table[14][1] = 0;
assign binom_table[14][2] = 0;
assign binom_table[14][3] = 0;
assign binom_table[14][4] = 0;
assign binom_table[14][5] = 0;
assign binom_table[14][6] = 0;
assign binom_table[14][7] = 0;
assign binom_table[14][8] = 0;
assign binom_table[14][9] = 0;
assign binom_table[14][10] = 0;
assign binom_table[14][11] = 0;
assign binom_table[14][12] = 0;
assign binom_table[14][13] = 0;
assign binom_table[14][14] = 1;
assign binom_table[14][15] = 15;
assign binom_table[14][16] = 120;
assign binom_table[14][17] = 680;
assign binom_table[14][18] = 3060;
assign binom_table[14][19] = 11628;
assign binom_table[14][20] = 38760;
assign binom_table[14][21] = 116280;
assign binom_table[14][22] = 319770;
assign binom_table[14][23] = 817190;
assign binom_table[14][24] = 1961256;
assign binom_table[14][25] = 4457400;
assign binom_table[14][26] = 9657700;
assign binom_table[14][27] = 20058300;
assign binom_table[14][28] = 40116600;
assign binom_table[14][29] = 77558760;
assign binom_table[14][30] = 145422675;
assign binom_table[14][31] = 265182525;
assign binom_table[14][32] = 471435600;

assign binom_table[15][1] = 0;
assign binom_table[15][2] = 0;
assign binom_table[15][3] = 0;
assign binom_table[15][4] = 0;
assign binom_table[15][5] = 0;
assign binom_table[15][6] = 0;
assign binom_table[15][7] = 0;
assign binom_table[15][8] = 0;
assign binom_table[15][9] = 0;
assign binom_table[15][10] = 0;
assign binom_table[15][11] = 0;
assign binom_table[15][12] = 0;
assign binom_table[15][13] = 0;
assign binom_table[15][14] = 0;
assign binom_table[15][15] = 1;
assign binom_table[15][16] = 16;
assign binom_table[15][17] = 136;
assign binom_table[15][18] = 816;
assign binom_table[15][19] = 3876;
assign binom_table[15][20] = 15504;
assign binom_table[15][21] = 54264;
assign binom_table[15][22] = 170544;
assign binom_table[15][23] = 490314;
assign binom_table[15][24] = 1307504;
assign binom_table[15][25] = 3268760;
assign binom_table[15][26] = 7726160;
assign binom_table[15][27] = 17383860;
assign binom_table[15][28] = 37442160;
assign binom_table[15][29] = 77558760;
assign binom_table[15][30] = 155117520;
assign binom_table[15][31] = 300540195;
assign binom_table[15][32] = 565722720;

assign binom_table[16][1] = 0;
assign binom_table[16][2] = 0;
assign binom_table[16][3] = 0;
assign binom_table[16][4] = 0;
assign binom_table[16][5] = 0;
assign binom_table[16][6] = 0;
assign binom_table[16][7] = 0;
assign binom_table[16][8] = 0;
assign binom_table[16][9] = 0;
assign binom_table[16][10] = 0;
assign binom_table[16][11] = 0;
assign binom_table[16][12] = 0;
assign binom_table[16][13] = 0;
assign binom_table[16][14] = 0;
assign binom_table[16][15] = 0;
assign binom_table[16][16] = 1;
assign binom_table[16][17] = 17;
assign binom_table[16][18] = 153;
assign binom_table[16][19] = 969;
assign binom_table[16][20] = 4845;
assign binom_table[16][21] = 20349;
assign binom_table[16][22] = 74613;
assign binom_table[16][23] = 245157;
assign binom_table[16][24] = 735471;
assign binom_table[16][25] = 2042975;
assign binom_table[16][26] = 5311735;
assign binom_table[16][27] = 13037895;
assign binom_table[16][28] = 30421755;
assign binom_table[16][29] = 67863915;
assign binom_table[16][30] = 145422675;
assign binom_table[16][31] = 300540195;
assign binom_table[16][32] = 601080390;

assign binom_table[17][1] = 0;
assign binom_table[17][2] = 0;
assign binom_table[17][3] = 0;
assign binom_table[17][4] = 0;
assign binom_table[17][5] = 0;
assign binom_table[17][6] = 0;
assign binom_table[17][7] = 0;
assign binom_table[17][8] = 0;
assign binom_table[17][9] = 0;
assign binom_table[17][10] = 0;
assign binom_table[17][11] = 0;
assign binom_table[17][12] = 0;
assign binom_table[17][13] = 0;
assign binom_table[17][14] = 0;
assign binom_table[17][15] = 0;
assign binom_table[17][16] = 0;
assign binom_table[17][17] = 1;
assign binom_table[17][18] = 18;
assign binom_table[17][19] = 171;
assign binom_table[17][20] = 1140;
assign binom_table[17][21] = 5985;
assign binom_table[17][22] = 26334;
assign binom_table[17][23] = 100947;
assign binom_table[17][24] = 346104;
assign binom_table[17][25] = 1081575;
assign binom_table[17][26] = 3124550;
assign binom_table[17][27] = 8436285;
assign binom_table[17][28] = 21474180;
assign binom_table[17][29] = 51895935;
assign binom_table[17][30] = 119759850;
assign binom_table[17][31] = 265182525;
assign binom_table[17][32] = 565722720;

assign binom_table[18][1] = 0;
assign binom_table[18][2] = 0;
assign binom_table[18][3] = 0;
assign binom_table[18][4] = 0;
assign binom_table[18][5] = 0;
assign binom_table[18][6] = 0;
assign binom_table[18][7] = 0;
assign binom_table[18][8] = 0;
assign binom_table[18][9] = 0;
assign binom_table[18][10] = 0;
assign binom_table[18][11] = 0;
assign binom_table[18][12] = 0;
assign binom_table[18][13] = 0;
assign binom_table[18][14] = 0;
assign binom_table[18][15] = 0;
assign binom_table[18][16] = 0;
assign binom_table[18][17] = 0;
assign binom_table[18][18] = 1;
assign binom_table[18][19] = 19;
assign binom_table[18][20] = 190;
assign binom_table[18][21] = 1330;
assign binom_table[18][22] = 7315;
assign binom_table[18][23] = 33649;
assign binom_table[18][24] = 134596;
assign binom_table[18][25] = 480700;
assign binom_table[18][26] = 1562275;
assign binom_table[18][27] = 4686825;
assign binom_table[18][28] = 13123110;
assign binom_table[18][29] = 34597290;
assign binom_table[18][30] = 86493225;
assign binom_table[18][31] = 206253075;
assign binom_table[18][32] = 471435600;

assign binom_table[19][1] = 0;
assign binom_table[19][2] = 0;
assign binom_table[19][3] = 0;
assign binom_table[19][4] = 0;
assign binom_table[19][5] = 0;
assign binom_table[19][6] = 0;
assign binom_table[19][7] = 0;
assign binom_table[19][8] = 0;
assign binom_table[19][9] = 0;
assign binom_table[19][10] = 0;
assign binom_table[19][11] = 0;
assign binom_table[19][12] = 0;
assign binom_table[19][13] = 0;
assign binom_table[19][14] = 0;
assign binom_table[19][15] = 0;
assign binom_table[19][16] = 0;
assign binom_table[19][17] = 0;
assign binom_table[19][18] = 0;
assign binom_table[19][19] = 1;
assign binom_table[19][20] = 20;
assign binom_table[19][21] = 210;
assign binom_table[19][22] = 1540;
assign binom_table[19][23] = 8855;
assign binom_table[19][24] = 42504;
assign binom_table[19][25] = 177100;
assign binom_table[19][26] = 657800;
assign binom_table[19][27] = 2220075;
assign binom_table[19][28] = 6906900;
assign binom_table[19][29] = 20030010;
assign binom_table[19][30] = 54627300;
assign binom_table[19][31] = 141120525;
assign binom_table[19][32] = 347373600;

assign binom_table[20][1] = 0;
assign binom_table[20][2] = 0;
assign binom_table[20][3] = 0;
assign binom_table[20][4] = 0;
assign binom_table[20][5] = 0;
assign binom_table[20][6] = 0;
assign binom_table[20][7] = 0;
assign binom_table[20][8] = 0;
assign binom_table[20][9] = 0;
assign binom_table[20][10] = 0;
assign binom_table[20][11] = 0;
assign binom_table[20][12] = 0;
assign binom_table[20][13] = 0;
assign binom_table[20][14] = 0;
assign binom_table[20][15] = 0;
assign binom_table[20][16] = 0;
assign binom_table[20][17] = 0;
assign binom_table[20][18] = 0;
assign binom_table[20][19] = 0;
assign binom_table[20][20] = 1;
assign binom_table[20][21] = 21;
assign binom_table[20][22] = 231;
assign binom_table[20][23] = 1771;
assign binom_table[20][24] = 10626;
assign binom_table[20][25] = 53130;
assign binom_table[20][26] = 230230;
assign binom_table[20][27] = 888030;
assign binom_table[20][28] = 3108105;
assign binom_table[20][29] = 10015005;
assign binom_table[20][30] = 30045015;
assign binom_table[20][31] = 84672315;
assign binom_table[20][32] = 225792840;

assign binom_table[21][1] = 0;
assign binom_table[21][2] = 0;
assign binom_table[21][3] = 0;
assign binom_table[21][4] = 0;
assign binom_table[21][5] = 0;
assign binom_table[21][6] = 0;
assign binom_table[21][7] = 0;
assign binom_table[21][8] = 0;
assign binom_table[21][9] = 0;
assign binom_table[21][10] = 0;
assign binom_table[21][11] = 0;
assign binom_table[21][12] = 0;
assign binom_table[21][13] = 0;
assign binom_table[21][14] = 0;
assign binom_table[21][15] = 0;
assign binom_table[21][16] = 0;
assign binom_table[21][17] = 0;
assign binom_table[21][18] = 0;
assign binom_table[21][19] = 0;
assign binom_table[21][20] = 0;
assign binom_table[21][21] = 1;
assign binom_table[21][22] = 22;
assign binom_table[21][23] = 253;
assign binom_table[21][24] = 2024;
assign binom_table[21][25] = 12650;
assign binom_table[21][26] = 65780;
assign binom_table[21][27] = 296010;
assign binom_table[21][28] = 1184040;
assign binom_table[21][29] = 4292145;
assign binom_table[21][30] = 14307150;
assign binom_table[21][31] = 44352165;
assign binom_table[21][32] = 129024480;

assign binom_table[22][1] = 0;
assign binom_table[22][2] = 0;
assign binom_table[22][3] = 0;
assign binom_table[22][4] = 0;
assign binom_table[22][5] = 0;
assign binom_table[22][6] = 0;
assign binom_table[22][7] = 0;
assign binom_table[22][8] = 0;
assign binom_table[22][9] = 0;
assign binom_table[22][10] = 0;
assign binom_table[22][11] = 0;
assign binom_table[22][12] = 0;
assign binom_table[22][13] = 0;
assign binom_table[22][14] = 0;
assign binom_table[22][15] = 0;
assign binom_table[22][16] = 0;
assign binom_table[22][17] = 0;
assign binom_table[22][18] = 0;
assign binom_table[22][19] = 0;
assign binom_table[22][20] = 0;
assign binom_table[22][21] = 0;
assign binom_table[22][22] = 1;
assign binom_table[22][23] = 23;
assign binom_table[22][24] = 276;
assign binom_table[22][25] = 2300;
assign binom_table[22][26] = 14950;
assign binom_table[22][27] = 80730;
assign binom_table[22][28] = 376740;
assign binom_table[22][29] = 1560780;
assign binom_table[22][30] = 5852925;
assign binom_table[22][31] = 20160075;
assign binom_table[22][32] = 64512240;

assign binom_table[23][1] = 0;
assign binom_table[23][2] = 0;
assign binom_table[23][3] = 0;
assign binom_table[23][4] = 0;
assign binom_table[23][5] = 0;
assign binom_table[23][6] = 0;
assign binom_table[23][7] = 0;
assign binom_table[23][8] = 0;
assign binom_table[23][9] = 0;
assign binom_table[23][10] = 0;
assign binom_table[23][11] = 0;
assign binom_table[23][12] = 0;
assign binom_table[23][13] = 0;
assign binom_table[23][14] = 0;
assign binom_table[23][15] = 0;
assign binom_table[23][16] = 0;
assign binom_table[23][17] = 0;
assign binom_table[23][18] = 0;
assign binom_table[23][19] = 0;
assign binom_table[23][20] = 0;
assign binom_table[23][21] = 0;
assign binom_table[23][22] = 0;
assign binom_table[23][23] = 1;
assign binom_table[23][24] = 24;
assign binom_table[23][25] = 300;
assign binom_table[23][26] = 2600;
assign binom_table[23][27] = 17550;
assign binom_table[23][28] = 98280;
assign binom_table[23][29] = 475020;
assign binom_table[23][30] = 2035800;
assign binom_table[23][31] = 7888725;
assign binom_table[23][32] = 28048800;

assign binom_table[24][1] = 0;
assign binom_table[24][2] = 0;
assign binom_table[24][3] = 0;
assign binom_table[24][4] = 0;
assign binom_table[24][5] = 0;
assign binom_table[24][6] = 0;
assign binom_table[24][7] = 0;
assign binom_table[24][8] = 0;
assign binom_table[24][9] = 0;
assign binom_table[24][10] = 0;
assign binom_table[24][11] = 0;
assign binom_table[24][12] = 0;
assign binom_table[24][13] = 0;
assign binom_table[24][14] = 0;
assign binom_table[24][15] = 0;
assign binom_table[24][16] = 0;
assign binom_table[24][17] = 0;
assign binom_table[24][18] = 0;
assign binom_table[24][19] = 0;
assign binom_table[24][20] = 0;
assign binom_table[24][21] = 0;
assign binom_table[24][22] = 0;
assign binom_table[24][23] = 0;
assign binom_table[24][24] = 1;
assign binom_table[24][25] = 25;
assign binom_table[24][26] = 325;
assign binom_table[24][27] = 2925;
assign binom_table[24][28] = 20475;
assign binom_table[24][29] = 118755;
assign binom_table[24][30] = 593775;
assign binom_table[24][31] = 2629575;
assign binom_table[24][32] = 10518300;

assign binom_table[25][1] = 0;
assign binom_table[25][2] = 0;
assign binom_table[25][3] = 0;
assign binom_table[25][4] = 0;
assign binom_table[25][5] = 0;
assign binom_table[25][6] = 0;
assign binom_table[25][7] = 0;
assign binom_table[25][8] = 0;
assign binom_table[25][9] = 0;
assign binom_table[25][10] = 0;
assign binom_table[25][11] = 0;
assign binom_table[25][12] = 0;
assign binom_table[25][13] = 0;
assign binom_table[25][14] = 0;
assign binom_table[25][15] = 0;
assign binom_table[25][16] = 0;
assign binom_table[25][17] = 0;
assign binom_table[25][18] = 0;
assign binom_table[25][19] = 0;
assign binom_table[25][20] = 0;
assign binom_table[25][21] = 0;
assign binom_table[25][22] = 0;
assign binom_table[25][23] = 0;
assign binom_table[25][24] = 0;
assign binom_table[25][25] = 1;
assign binom_table[25][26] = 26;
assign binom_table[25][27] = 351;
assign binom_table[25][28] = 3276;
assign binom_table[25][29] = 23751;
assign binom_table[25][30] = 142506;
assign binom_table[25][31] = 736281;
assign binom_table[25][32] = 3365856;

assign binom_table[26][1] = 0;
assign binom_table[26][2] = 0;
assign binom_table[26][3] = 0;
assign binom_table[26][4] = 0;
assign binom_table[26][5] = 0;
assign binom_table[26][6] = 0;
assign binom_table[26][7] = 0;
assign binom_table[26][8] = 0;
assign binom_table[26][9] = 0;
assign binom_table[26][10] = 0;
assign binom_table[26][11] = 0;
assign binom_table[26][12] = 0;
assign binom_table[26][13] = 0;
assign binom_table[26][14] = 0;
assign binom_table[26][15] = 0;
assign binom_table[26][16] = 0;
assign binom_table[26][17] = 0;
assign binom_table[26][18] = 0;
assign binom_table[26][19] = 0;
assign binom_table[26][20] = 0;
assign binom_table[26][21] = 0;
assign binom_table[26][22] = 0;
assign binom_table[26][23] = 0;
assign binom_table[26][24] = 0;
assign binom_table[26][25] = 0;
assign binom_table[26][26] = 1;
assign binom_table[26][27] = 27;
assign binom_table[26][28] = 378;
assign binom_table[26][29] = 3654;
assign binom_table[26][30] = 27405;
assign binom_table[26][31] = 169911;
assign binom_table[26][32] = 906192;

assign binom_table[27][1] = 0;
assign binom_table[27][2] = 0;
assign binom_table[27][3] = 0;
assign binom_table[27][4] = 0;
assign binom_table[27][5] = 0;
assign binom_table[27][6] = 0;
assign binom_table[27][7] = 0;
assign binom_table[27][8] = 0;
assign binom_table[27][9] = 0;
assign binom_table[27][10] = 0;
assign binom_table[27][11] = 0;
assign binom_table[27][12] = 0;
assign binom_table[27][13] = 0;
assign binom_table[27][14] = 0;
assign binom_table[27][15] = 0;
assign binom_table[27][16] = 0;
assign binom_table[27][17] = 0;
assign binom_table[27][18] = 0;
assign binom_table[27][19] = 0;
assign binom_table[27][20] = 0;
assign binom_table[27][21] = 0;
assign binom_table[27][22] = 0;
assign binom_table[27][23] = 0;
assign binom_table[27][24] = 0;
assign binom_table[27][25] = 0;
assign binom_table[27][26] = 0;
assign binom_table[27][27] = 1;
assign binom_table[27][28] = 28;
assign binom_table[27][29] = 406;
assign binom_table[27][30] = 4060;
assign binom_table[27][31] = 31465;
assign binom_table[27][32] = 201376;

assign binom_table[28][1] = 0;
assign binom_table[28][2] = 0;
assign binom_table[28][3] = 0;
assign binom_table[28][4] = 0;
assign binom_table[28][5] = 0;
assign binom_table[28][6] = 0;
assign binom_table[28][7] = 0;
assign binom_table[28][8] = 0;
assign binom_table[28][9] = 0;
assign binom_table[28][10] = 0;
assign binom_table[28][11] = 0;
assign binom_table[28][12] = 0;
assign binom_table[28][13] = 0;
assign binom_table[28][14] = 0;
assign binom_table[28][15] = 0;
assign binom_table[28][16] = 0;
assign binom_table[28][17] = 0;
assign binom_table[28][18] = 0;
assign binom_table[28][19] = 0;
assign binom_table[28][20] = 0;
assign binom_table[28][21] = 0;
assign binom_table[28][22] = 0;
assign binom_table[28][23] = 0;
assign binom_table[28][24] = 0;
assign binom_table[28][25] = 0;
assign binom_table[28][26] = 0;
assign binom_table[28][27] = 0;
assign binom_table[28][28] = 1;
assign binom_table[28][29] = 29;
assign binom_table[28][30] = 435;
assign binom_table[28][31] = 4495;
assign binom_table[28][32] = 35960;

assign binom_table[29][1] = 0;
assign binom_table[29][2] = 0;
assign binom_table[29][3] = 0;
assign binom_table[29][4] = 0;
assign binom_table[29][5] = 0;
assign binom_table[29][6] = 0;
assign binom_table[29][7] = 0;
assign binom_table[29][8] = 0;
assign binom_table[29][9] = 0;
assign binom_table[29][10] = 0;
assign binom_table[29][11] = 0;
assign binom_table[29][12] = 0;
assign binom_table[29][13] = 0;
assign binom_table[29][14] = 0;
assign binom_table[29][15] = 0;
assign binom_table[29][16] = 0;
assign binom_table[29][17] = 0;
assign binom_table[29][18] = 0;
assign binom_table[29][19] = 0;
assign binom_table[29][20] = 0;
assign binom_table[29][21] = 0;
assign binom_table[29][22] = 0;
assign binom_table[29][23] = 0;
assign binom_table[29][24] = 0;
assign binom_table[29][25] = 0;
assign binom_table[29][26] = 0;
assign binom_table[29][27] = 0;
assign binom_table[29][28] = 0;
assign binom_table[29][29] = 1;
assign binom_table[29][30] = 30;
assign binom_table[29][31] = 465;
assign binom_table[29][32] = 4960;

assign binom_table[30][1] = 0;
assign binom_table[30][2] = 0;
assign binom_table[30][3] = 0;
assign binom_table[30][4] = 0;
assign binom_table[30][5] = 0;
assign binom_table[30][6] = 0;
assign binom_table[30][7] = 0;
assign binom_table[30][8] = 0;
assign binom_table[30][9] = 0;
assign binom_table[30][10] = 0;
assign binom_table[30][11] = 0;
assign binom_table[30][12] = 0;
assign binom_table[30][13] = 0;
assign binom_table[30][14] = 0;
assign binom_table[30][15] = 0;
assign binom_table[30][16] = 0;
assign binom_table[30][17] = 0;
assign binom_table[30][18] = 0;
assign binom_table[30][19] = 0;
assign binom_table[30][20] = 0;
assign binom_table[30][21] = 0;
assign binom_table[30][22] = 0;
assign binom_table[30][23] = 0;
assign binom_table[30][24] = 0;
assign binom_table[30][25] = 0;
assign binom_table[30][26] = 0;
assign binom_table[30][27] = 0;
assign binom_table[30][28] = 0;
assign binom_table[30][29] = 0;
assign binom_table[30][30] = 1;
assign binom_table[30][31] = 31;
assign binom_table[30][32] = 496;

assign binom_table[31][1] = 0;
assign binom_table[31][2] = 0;
assign binom_table[31][3] = 0;
assign binom_table[31][4] = 0;
assign binom_table[31][5] = 0;
assign binom_table[31][6] = 0;
assign binom_table[31][7] = 0;
assign binom_table[31][8] = 0;
assign binom_table[31][9] = 0;
assign binom_table[31][10] = 0;
assign binom_table[31][11] = 0;
assign binom_table[31][12] = 0;
assign binom_table[31][13] = 0;
assign binom_table[31][14] = 0;
assign binom_table[31][15] = 0;
assign binom_table[31][16] = 0;
assign binom_table[31][17] = 0;
assign binom_table[31][18] = 0;
assign binom_table[31][19] = 0;
assign binom_table[31][20] = 0;
assign binom_table[31][21] = 0;
assign binom_table[31][22] = 0;
assign binom_table[31][23] = 0;
assign binom_table[31][24] = 0;
assign binom_table[31][25] = 0;
assign binom_table[31][26] = 0;
assign binom_table[31][27] = 0;
assign binom_table[31][28] = 0;
assign binom_table[31][29] = 0;
assign binom_table[31][30] = 0;
assign binom_table[31][31] = 1;
assign binom_table[31][32] = 32;

assign binom_table[32][1] = 0;
assign binom_table[32][2] = 0;
assign binom_table[32][3] = 0;
assign binom_table[32][4] = 0;
assign binom_table[32][5] = 0;
assign binom_table[32][6] = 0;
assign binom_table[32][7] = 0;
assign binom_table[32][8] = 0;
assign binom_table[32][9] = 0;
assign binom_table[32][10] = 0;
assign binom_table[32][11] = 0;
assign binom_table[32][12] = 0;
assign binom_table[32][13] = 0;
assign binom_table[32][14] = 0;
assign binom_table[32][15] = 0;
assign binom_table[32][16] = 0;
assign binom_table[32][17] = 0;
assign binom_table[32][18] = 0;
assign binom_table[32][19] = 0;
assign binom_table[32][20] = 0;
assign binom_table[32][21] = 0;
assign binom_table[32][22] = 0;
assign binom_table[32][23] = 0;
assign binom_table[32][24] = 0;
assign binom_table[32][25] = 0;
assign binom_table[32][26] = 0;
assign binom_table[32][27] = 0;
assign binom_table[32][28] = 0;
assign binom_table[32][29] = 0;
assign binom_table[32][30] = 0;
assign binom_table[32][31] = 0;
assign binom_table[32][32] = 1;

assign bits[1][1] = num > binom_table[1][1];
assign bits[1][2] = num > binom_table[1][2];
assign bits[1][3] = num > binom_table[1][3];
assign bits[1][4] = num > binom_table[1][4];
assign bits[1][5] = num > binom_table[1][5];
assign bits[1][6] = num > binom_table[1][6];
assign bits[1][7] = num > binom_table[1][7];
assign bits[1][8] = num > binom_table[1][8];
assign bits[1][9] = num > binom_table[1][9];
assign bits[1][10] = num > binom_table[1][10];
assign bits[1][11] = num > binom_table[1][11];
assign bits[1][12] = num > binom_table[1][12];
assign bits[1][13] = num > binom_table[1][13];
assign bits[1][14] = num > binom_table[1][14];
assign bits[1][15] = num > binom_table[1][15];
assign bits[1][16] = num > binom_table[1][16];
assign bits[1][17] = num > binom_table[1][17];
assign bits[1][18] = num > binom_table[1][18];
assign bits[1][19] = num > binom_table[1][19];
assign bits[1][20] = num > binom_table[1][20];
assign bits[1][21] = num > binom_table[1][21];
assign bits[1][22] = num > binom_table[1][22];
assign bits[1][23] = num > binom_table[1][23];
assign bits[1][24] = num > binom_table[1][24];
assign bits[1][25] = num > binom_table[1][25];
assign bits[1][26] = num > binom_table[1][26];
assign bits[1][27] = num > binom_table[1][27];
assign bits[1][28] = num > binom_table[1][28];
assign bits[1][29] = num > binom_table[1][29];
assign bits[1][30] = num > binom_table[1][30];
assign bits[1][31] = num > binom_table[1][31];
assign bits[1][32] = num > binom_table[1][32];

assign bits[2][1] = num > binom_table[2][1];
assign bits[2][2] = num > binom_table[2][2];
assign bits[2][3] = num > binom_table[2][3];
assign bits[2][4] = num > binom_table[2][4];
assign bits[2][5] = num > binom_table[2][5];
assign bits[2][6] = num > binom_table[2][6];
assign bits[2][7] = num > binom_table[2][7];
assign bits[2][8] = num > binom_table[2][8];
assign bits[2][9] = num > binom_table[2][9];
assign bits[2][10] = num > binom_table[2][10];
assign bits[2][11] = num > binom_table[2][11];
assign bits[2][12] = num > binom_table[2][12];
assign bits[2][13] = num > binom_table[2][13];
assign bits[2][14] = num > binom_table[2][14];
assign bits[2][15] = num > binom_table[2][15];
assign bits[2][16] = num > binom_table[2][16];
assign bits[2][17] = num > binom_table[2][17];
assign bits[2][18] = num > binom_table[2][18];
assign bits[2][19] = num > binom_table[2][19];
assign bits[2][20] = num > binom_table[2][20];
assign bits[2][21] = num > binom_table[2][21];
assign bits[2][22] = num > binom_table[2][22];
assign bits[2][23] = num > binom_table[2][23];
assign bits[2][24] = num > binom_table[2][24];
assign bits[2][25] = num > binom_table[2][25];
assign bits[2][26] = num > binom_table[2][26];
assign bits[2][27] = num > binom_table[2][27];
assign bits[2][28] = num > binom_table[2][28];
assign bits[2][29] = num > binom_table[2][29];
assign bits[2][30] = num > binom_table[2][30];
assign bits[2][31] = num > binom_table[2][31];
assign bits[2][32] = num > binom_table[2][32];

assign bits[3][1] = num > binom_table[3][1];
assign bits[3][2] = num > binom_table[3][2];
assign bits[3][3] = num > binom_table[3][3];
assign bits[3][4] = num > binom_table[3][4];
assign bits[3][5] = num > binom_table[3][5];
assign bits[3][6] = num > binom_table[3][6];
assign bits[3][7] = num > binom_table[3][7];
assign bits[3][8] = num > binom_table[3][8];
assign bits[3][9] = num > binom_table[3][9];
assign bits[3][10] = num > binom_table[3][10];
assign bits[3][11] = num > binom_table[3][11];
assign bits[3][12] = num > binom_table[3][12];
assign bits[3][13] = num > binom_table[3][13];
assign bits[3][14] = num > binom_table[3][14];
assign bits[3][15] = num > binom_table[3][15];
assign bits[3][16] = num > binom_table[3][16];
assign bits[3][17] = num > binom_table[3][17];
assign bits[3][18] = num > binom_table[3][18];
assign bits[3][19] = num > binom_table[3][19];
assign bits[3][20] = num > binom_table[3][20];
assign bits[3][21] = num > binom_table[3][21];
assign bits[3][22] = num > binom_table[3][22];
assign bits[3][23] = num > binom_table[3][23];
assign bits[3][24] = num > binom_table[3][24];
assign bits[3][25] = num > binom_table[3][25];
assign bits[3][26] = num > binom_table[3][26];
assign bits[3][27] = num > binom_table[3][27];
assign bits[3][28] = num > binom_table[3][28];
assign bits[3][29] = num > binom_table[3][29];
assign bits[3][30] = num > binom_table[3][30];
assign bits[3][31] = num > binom_table[3][31];
assign bits[3][32] = num > binom_table[3][32];

assign bits[4][1] = num > binom_table[4][1];
assign bits[4][2] = num > binom_table[4][2];
assign bits[4][3] = num > binom_table[4][3];
assign bits[4][4] = num > binom_table[4][4];
assign bits[4][5] = num > binom_table[4][5];
assign bits[4][6] = num > binom_table[4][6];
assign bits[4][7] = num > binom_table[4][7];
assign bits[4][8] = num > binom_table[4][8];
assign bits[4][9] = num > binom_table[4][9];
assign bits[4][10] = num > binom_table[4][10];
assign bits[4][11] = num > binom_table[4][11];
assign bits[4][12] = num > binom_table[4][12];
assign bits[4][13] = num > binom_table[4][13];
assign bits[4][14] = num > binom_table[4][14];
assign bits[4][15] = num > binom_table[4][15];
assign bits[4][16] = num > binom_table[4][16];
assign bits[4][17] = num > binom_table[4][17];
assign bits[4][18] = num > binom_table[4][18];
assign bits[4][19] = num > binom_table[4][19];
assign bits[4][20] = num > binom_table[4][20];
assign bits[4][21] = num > binom_table[4][21];
assign bits[4][22] = num > binom_table[4][22];
assign bits[4][23] = num > binom_table[4][23];
assign bits[4][24] = num > binom_table[4][24];
assign bits[4][25] = num > binom_table[4][25];
assign bits[4][26] = num > binom_table[4][26];
assign bits[4][27] = num > binom_table[4][27];
assign bits[4][28] = num > binom_table[4][28];
assign bits[4][29] = num > binom_table[4][29];
assign bits[4][30] = num > binom_table[4][30];
assign bits[4][31] = num > binom_table[4][31];
assign bits[4][32] = num > binom_table[4][32];

assign bits[5][1] = num > binom_table[5][1];
assign bits[5][2] = num > binom_table[5][2];
assign bits[5][3] = num > binom_table[5][3];
assign bits[5][4] = num > binom_table[5][4];
assign bits[5][5] = num > binom_table[5][5];
assign bits[5][6] = num > binom_table[5][6];
assign bits[5][7] = num > binom_table[5][7];
assign bits[5][8] = num > binom_table[5][8];
assign bits[5][9] = num > binom_table[5][9];
assign bits[5][10] = num > binom_table[5][10];
assign bits[5][11] = num > binom_table[5][11];
assign bits[5][12] = num > binom_table[5][12];
assign bits[5][13] = num > binom_table[5][13];
assign bits[5][14] = num > binom_table[5][14];
assign bits[5][15] = num > binom_table[5][15];
assign bits[5][16] = num > binom_table[5][16];
assign bits[5][17] = num > binom_table[5][17];
assign bits[5][18] = num > binom_table[5][18];
assign bits[5][19] = num > binom_table[5][19];
assign bits[5][20] = num > binom_table[5][20];
assign bits[5][21] = num > binom_table[5][21];
assign bits[5][22] = num > binom_table[5][22];
assign bits[5][23] = num > binom_table[5][23];
assign bits[5][24] = num > binom_table[5][24];
assign bits[5][25] = num > binom_table[5][25];
assign bits[5][26] = num > binom_table[5][26];
assign bits[5][27] = num > binom_table[5][27];
assign bits[5][28] = num > binom_table[5][28];
assign bits[5][29] = num > binom_table[5][29];
assign bits[5][30] = num > binom_table[5][30];
assign bits[5][31] = num > binom_table[5][31];
assign bits[5][32] = num > binom_table[5][32];

assign bits[6][1] = num > binom_table[6][1];
assign bits[6][2] = num > binom_table[6][2];
assign bits[6][3] = num > binom_table[6][3];
assign bits[6][4] = num > binom_table[6][4];
assign bits[6][5] = num > binom_table[6][5];
assign bits[6][6] = num > binom_table[6][6];
assign bits[6][7] = num > binom_table[6][7];
assign bits[6][8] = num > binom_table[6][8];
assign bits[6][9] = num > binom_table[6][9];
assign bits[6][10] = num > binom_table[6][10];
assign bits[6][11] = num > binom_table[6][11];
assign bits[6][12] = num > binom_table[6][12];
assign bits[6][13] = num > binom_table[6][13];
assign bits[6][14] = num > binom_table[6][14];
assign bits[6][15] = num > binom_table[6][15];
assign bits[6][16] = num > binom_table[6][16];
assign bits[6][17] = num > binom_table[6][17];
assign bits[6][18] = num > binom_table[6][18];
assign bits[6][19] = num > binom_table[6][19];
assign bits[6][20] = num > binom_table[6][20];
assign bits[6][21] = num > binom_table[6][21];
assign bits[6][22] = num > binom_table[6][22];
assign bits[6][23] = num > binom_table[6][23];
assign bits[6][24] = num > binom_table[6][24];
assign bits[6][25] = num > binom_table[6][25];
assign bits[6][26] = num > binom_table[6][26];
assign bits[6][27] = num > binom_table[6][27];
assign bits[6][28] = num > binom_table[6][28];
assign bits[6][29] = num > binom_table[6][29];
assign bits[6][30] = num > binom_table[6][30];
assign bits[6][31] = num > binom_table[6][31];
assign bits[6][32] = num > binom_table[6][32];

assign bits[7][1] = num > binom_table[7][1];
assign bits[7][2] = num > binom_table[7][2];
assign bits[7][3] = num > binom_table[7][3];
assign bits[7][4] = num > binom_table[7][4];
assign bits[7][5] = num > binom_table[7][5];
assign bits[7][6] = num > binom_table[7][6];
assign bits[7][7] = num > binom_table[7][7];
assign bits[7][8] = num > binom_table[7][8];
assign bits[7][9] = num > binom_table[7][9];
assign bits[7][10] = num > binom_table[7][10];
assign bits[7][11] = num > binom_table[7][11];
assign bits[7][12] = num > binom_table[7][12];
assign bits[7][13] = num > binom_table[7][13];
assign bits[7][14] = num > binom_table[7][14];
assign bits[7][15] = num > binom_table[7][15];
assign bits[7][16] = num > binom_table[7][16];
assign bits[7][17] = num > binom_table[7][17];
assign bits[7][18] = num > binom_table[7][18];
assign bits[7][19] = num > binom_table[7][19];
assign bits[7][20] = num > binom_table[7][20];
assign bits[7][21] = num > binom_table[7][21];
assign bits[7][22] = num > binom_table[7][22];
assign bits[7][23] = num > binom_table[7][23];
assign bits[7][24] = num > binom_table[7][24];
assign bits[7][25] = num > binom_table[7][25];
assign bits[7][26] = num > binom_table[7][26];
assign bits[7][27] = num > binom_table[7][27];
assign bits[7][28] = num > binom_table[7][28];
assign bits[7][29] = num > binom_table[7][29];
assign bits[7][30] = num > binom_table[7][30];
assign bits[7][31] = num > binom_table[7][31];
assign bits[7][32] = num > binom_table[7][32];

assign bits[8][1] = num > binom_table[8][1];
assign bits[8][2] = num > binom_table[8][2];
assign bits[8][3] = num > binom_table[8][3];
assign bits[8][4] = num > binom_table[8][4];
assign bits[8][5] = num > binom_table[8][5];
assign bits[8][6] = num > binom_table[8][6];
assign bits[8][7] = num > binom_table[8][7];
assign bits[8][8] = num > binom_table[8][8];
assign bits[8][9] = num > binom_table[8][9];
assign bits[8][10] = num > binom_table[8][10];
assign bits[8][11] = num > binom_table[8][11];
assign bits[8][12] = num > binom_table[8][12];
assign bits[8][13] = num > binom_table[8][13];
assign bits[8][14] = num > binom_table[8][14];
assign bits[8][15] = num > binom_table[8][15];
assign bits[8][16] = num > binom_table[8][16];
assign bits[8][17] = num > binom_table[8][17];
assign bits[8][18] = num > binom_table[8][18];
assign bits[8][19] = num > binom_table[8][19];
assign bits[8][20] = num > binom_table[8][20];
assign bits[8][21] = num > binom_table[8][21];
assign bits[8][22] = num > binom_table[8][22];
assign bits[8][23] = num > binom_table[8][23];
assign bits[8][24] = num > binom_table[8][24];
assign bits[8][25] = num > binom_table[8][25];
assign bits[8][26] = num > binom_table[8][26];
assign bits[8][27] = num > binom_table[8][27];
assign bits[8][28] = num > binom_table[8][28];
assign bits[8][29] = num > binom_table[8][29];
assign bits[8][30] = num > binom_table[8][30];
assign bits[8][31] = num > binom_table[8][31];
assign bits[8][32] = num > binom_table[8][32];

assign bits[9][1] = num > binom_table[9][1];
assign bits[9][2] = num > binom_table[9][2];
assign bits[9][3] = num > binom_table[9][3];
assign bits[9][4] = num > binom_table[9][4];
assign bits[9][5] = num > binom_table[9][5];
assign bits[9][6] = num > binom_table[9][6];
assign bits[9][7] = num > binom_table[9][7];
assign bits[9][8] = num > binom_table[9][8];
assign bits[9][9] = num > binom_table[9][9];
assign bits[9][10] = num > binom_table[9][10];
assign bits[9][11] = num > binom_table[9][11];
assign bits[9][12] = num > binom_table[9][12];
assign bits[9][13] = num > binom_table[9][13];
assign bits[9][14] = num > binom_table[9][14];
assign bits[9][15] = num > binom_table[9][15];
assign bits[9][16] = num > binom_table[9][16];
assign bits[9][17] = num > binom_table[9][17];
assign bits[9][18] = num > binom_table[9][18];
assign bits[9][19] = num > binom_table[9][19];
assign bits[9][20] = num > binom_table[9][20];
assign bits[9][21] = num > binom_table[9][21];
assign bits[9][22] = num > binom_table[9][22];
assign bits[9][23] = num > binom_table[9][23];
assign bits[9][24] = num > binom_table[9][24];
assign bits[9][25] = num > binom_table[9][25];
assign bits[9][26] = num > binom_table[9][26];
assign bits[9][27] = num > binom_table[9][27];
assign bits[9][28] = num > binom_table[9][28];
assign bits[9][29] = num > binom_table[9][29];
assign bits[9][30] = num > binom_table[9][30];
assign bits[9][31] = num > binom_table[9][31];
assign bits[9][32] = num > binom_table[9][32];

assign bits[10][1] = num > binom_table[10][1];
assign bits[10][2] = num > binom_table[10][2];
assign bits[10][3] = num > binom_table[10][3];
assign bits[10][4] = num > binom_table[10][4];
assign bits[10][5] = num > binom_table[10][5];
assign bits[10][6] = num > binom_table[10][6];
assign bits[10][7] = num > binom_table[10][7];
assign bits[10][8] = num > binom_table[10][8];
assign bits[10][9] = num > binom_table[10][9];
assign bits[10][10] = num > binom_table[10][10];
assign bits[10][11] = num > binom_table[10][11];
assign bits[10][12] = num > binom_table[10][12];
assign bits[10][13] = num > binom_table[10][13];
assign bits[10][14] = num > binom_table[10][14];
assign bits[10][15] = num > binom_table[10][15];
assign bits[10][16] = num > binom_table[10][16];
assign bits[10][17] = num > binom_table[10][17];
assign bits[10][18] = num > binom_table[10][18];
assign bits[10][19] = num > binom_table[10][19];
assign bits[10][20] = num > binom_table[10][20];
assign bits[10][21] = num > binom_table[10][21];
assign bits[10][22] = num > binom_table[10][22];
assign bits[10][23] = num > binom_table[10][23];
assign bits[10][24] = num > binom_table[10][24];
assign bits[10][25] = num > binom_table[10][25];
assign bits[10][26] = num > binom_table[10][26];
assign bits[10][27] = num > binom_table[10][27];
assign bits[10][28] = num > binom_table[10][28];
assign bits[10][29] = num > binom_table[10][29];
assign bits[10][30] = num > binom_table[10][30];
assign bits[10][31] = num > binom_table[10][31];
assign bits[10][32] = num > binom_table[10][32];

assign bits[11][1] = num > binom_table[11][1];
assign bits[11][2] = num > binom_table[11][2];
assign bits[11][3] = num > binom_table[11][3];
assign bits[11][4] = num > binom_table[11][4];
assign bits[11][5] = num > binom_table[11][5];
assign bits[11][6] = num > binom_table[11][6];
assign bits[11][7] = num > binom_table[11][7];
assign bits[11][8] = num > binom_table[11][8];
assign bits[11][9] = num > binom_table[11][9];
assign bits[11][10] = num > binom_table[11][10];
assign bits[11][11] = num > binom_table[11][11];
assign bits[11][12] = num > binom_table[11][12];
assign bits[11][13] = num > binom_table[11][13];
assign bits[11][14] = num > binom_table[11][14];
assign bits[11][15] = num > binom_table[11][15];
assign bits[11][16] = num > binom_table[11][16];
assign bits[11][17] = num > binom_table[11][17];
assign bits[11][18] = num > binom_table[11][18];
assign bits[11][19] = num > binom_table[11][19];
assign bits[11][20] = num > binom_table[11][20];
assign bits[11][21] = num > binom_table[11][21];
assign bits[11][22] = num > binom_table[11][22];
assign bits[11][23] = num > binom_table[11][23];
assign bits[11][24] = num > binom_table[11][24];
assign bits[11][25] = num > binom_table[11][25];
assign bits[11][26] = num > binom_table[11][26];
assign bits[11][27] = num > binom_table[11][27];
assign bits[11][28] = num > binom_table[11][28];
assign bits[11][29] = num > binom_table[11][29];
assign bits[11][30] = num > binom_table[11][30];
assign bits[11][31] = num > binom_table[11][31];
assign bits[11][32] = num > binom_table[11][32];

assign bits[12][1] = num > binom_table[12][1];
assign bits[12][2] = num > binom_table[12][2];
assign bits[12][3] = num > binom_table[12][3];
assign bits[12][4] = num > binom_table[12][4];
assign bits[12][5] = num > binom_table[12][5];
assign bits[12][6] = num > binom_table[12][6];
assign bits[12][7] = num > binom_table[12][7];
assign bits[12][8] = num > binom_table[12][8];
assign bits[12][9] = num > binom_table[12][9];
assign bits[12][10] = num > binom_table[12][10];
assign bits[12][11] = num > binom_table[12][11];
assign bits[12][12] = num > binom_table[12][12];
assign bits[12][13] = num > binom_table[12][13];
assign bits[12][14] = num > binom_table[12][14];
assign bits[12][15] = num > binom_table[12][15];
assign bits[12][16] = num > binom_table[12][16];
assign bits[12][17] = num > binom_table[12][17];
assign bits[12][18] = num > binom_table[12][18];
assign bits[12][19] = num > binom_table[12][19];
assign bits[12][20] = num > binom_table[12][20];
assign bits[12][21] = num > binom_table[12][21];
assign bits[12][22] = num > binom_table[12][22];
assign bits[12][23] = num > binom_table[12][23];
assign bits[12][24] = num > binom_table[12][24];
assign bits[12][25] = num > binom_table[12][25];
assign bits[12][26] = num > binom_table[12][26];
assign bits[12][27] = num > binom_table[12][27];
assign bits[12][28] = num > binom_table[12][28];
assign bits[12][29] = num > binom_table[12][29];
assign bits[12][30] = num > binom_table[12][30];
assign bits[12][31] = num > binom_table[12][31];
assign bits[12][32] = num > binom_table[12][32];

assign bits[13][1] = num > binom_table[13][1];
assign bits[13][2] = num > binom_table[13][2];
assign bits[13][3] = num > binom_table[13][3];
assign bits[13][4] = num > binom_table[13][4];
assign bits[13][5] = num > binom_table[13][5];
assign bits[13][6] = num > binom_table[13][6];
assign bits[13][7] = num > binom_table[13][7];
assign bits[13][8] = num > binom_table[13][8];
assign bits[13][9] = num > binom_table[13][9];
assign bits[13][10] = num > binom_table[13][10];
assign bits[13][11] = num > binom_table[13][11];
assign bits[13][12] = num > binom_table[13][12];
assign bits[13][13] = num > binom_table[13][13];
assign bits[13][14] = num > binom_table[13][14];
assign bits[13][15] = num > binom_table[13][15];
assign bits[13][16] = num > binom_table[13][16];
assign bits[13][17] = num > binom_table[13][17];
assign bits[13][18] = num > binom_table[13][18];
assign bits[13][19] = num > binom_table[13][19];
assign bits[13][20] = num > binom_table[13][20];
assign bits[13][21] = num > binom_table[13][21];
assign bits[13][22] = num > binom_table[13][22];
assign bits[13][23] = num > binom_table[13][23];
assign bits[13][24] = num > binom_table[13][24];
assign bits[13][25] = num > binom_table[13][25];
assign bits[13][26] = num > binom_table[13][26];
assign bits[13][27] = num > binom_table[13][27];
assign bits[13][28] = num > binom_table[13][28];
assign bits[13][29] = num > binom_table[13][29];
assign bits[13][30] = num > binom_table[13][30];
assign bits[13][31] = num > binom_table[13][31];
assign bits[13][32] = num > binom_table[13][32];

assign bits[14][1] = num > binom_table[14][1];
assign bits[14][2] = num > binom_table[14][2];
assign bits[14][3] = num > binom_table[14][3];
assign bits[14][4] = num > binom_table[14][4];
assign bits[14][5] = num > binom_table[14][5];
assign bits[14][6] = num > binom_table[14][6];
assign bits[14][7] = num > binom_table[14][7];
assign bits[14][8] = num > binom_table[14][8];
assign bits[14][9] = num > binom_table[14][9];
assign bits[14][10] = num > binom_table[14][10];
assign bits[14][11] = num > binom_table[14][11];
assign bits[14][12] = num > binom_table[14][12];
assign bits[14][13] = num > binom_table[14][13];
assign bits[14][14] = num > binom_table[14][14];
assign bits[14][15] = num > binom_table[14][15];
assign bits[14][16] = num > binom_table[14][16];
assign bits[14][17] = num > binom_table[14][17];
assign bits[14][18] = num > binom_table[14][18];
assign bits[14][19] = num > binom_table[14][19];
assign bits[14][20] = num > binom_table[14][20];
assign bits[14][21] = num > binom_table[14][21];
assign bits[14][22] = num > binom_table[14][22];
assign bits[14][23] = num > binom_table[14][23];
assign bits[14][24] = num > binom_table[14][24];
assign bits[14][25] = num > binom_table[14][25];
assign bits[14][26] = num > binom_table[14][26];
assign bits[14][27] = num > binom_table[14][27];
assign bits[14][28] = num > binom_table[14][28];
assign bits[14][29] = num > binom_table[14][29];
assign bits[14][30] = num > binom_table[14][30];
assign bits[14][31] = num > binom_table[14][31];
assign bits[14][32] = num > binom_table[14][32];

assign bits[15][1] = num > binom_table[15][1];
assign bits[15][2] = num > binom_table[15][2];
assign bits[15][3] = num > binom_table[15][3];
assign bits[15][4] = num > binom_table[15][4];
assign bits[15][5] = num > binom_table[15][5];
assign bits[15][6] = num > binom_table[15][6];
assign bits[15][7] = num > binom_table[15][7];
assign bits[15][8] = num > binom_table[15][8];
assign bits[15][9] = num > binom_table[15][9];
assign bits[15][10] = num > binom_table[15][10];
assign bits[15][11] = num > binom_table[15][11];
assign bits[15][12] = num > binom_table[15][12];
assign bits[15][13] = num > binom_table[15][13];
assign bits[15][14] = num > binom_table[15][14];
assign bits[15][15] = num > binom_table[15][15];
assign bits[15][16] = num > binom_table[15][16];
assign bits[15][17] = num > binom_table[15][17];
assign bits[15][18] = num > binom_table[15][18];
assign bits[15][19] = num > binom_table[15][19];
assign bits[15][20] = num > binom_table[15][20];
assign bits[15][21] = num > binom_table[15][21];
assign bits[15][22] = num > binom_table[15][22];
assign bits[15][23] = num > binom_table[15][23];
assign bits[15][24] = num > binom_table[15][24];
assign bits[15][25] = num > binom_table[15][25];
assign bits[15][26] = num > binom_table[15][26];
assign bits[15][27] = num > binom_table[15][27];
assign bits[15][28] = num > binom_table[15][28];
assign bits[15][29] = num > binom_table[15][29];
assign bits[15][30] = num > binom_table[15][30];
assign bits[15][31] = num > binom_table[15][31];
assign bits[15][32] = num > binom_table[15][32];

assign bits[16][1] = num > binom_table[16][1];
assign bits[16][2] = num > binom_table[16][2];
assign bits[16][3] = num > binom_table[16][3];
assign bits[16][4] = num > binom_table[16][4];
assign bits[16][5] = num > binom_table[16][5];
assign bits[16][6] = num > binom_table[16][6];
assign bits[16][7] = num > binom_table[16][7];
assign bits[16][8] = num > binom_table[16][8];
assign bits[16][9] = num > binom_table[16][9];
assign bits[16][10] = num > binom_table[16][10];
assign bits[16][11] = num > binom_table[16][11];
assign bits[16][12] = num > binom_table[16][12];
assign bits[16][13] = num > binom_table[16][13];
assign bits[16][14] = num > binom_table[16][14];
assign bits[16][15] = num > binom_table[16][15];
assign bits[16][16] = num > binom_table[16][16];
assign bits[16][17] = num > binom_table[16][17];
assign bits[16][18] = num > binom_table[16][18];
assign bits[16][19] = num > binom_table[16][19];
assign bits[16][20] = num > binom_table[16][20];
assign bits[16][21] = num > binom_table[16][21];
assign bits[16][22] = num > binom_table[16][22];
assign bits[16][23] = num > binom_table[16][23];
assign bits[16][24] = num > binom_table[16][24];
assign bits[16][25] = num > binom_table[16][25];
assign bits[16][26] = num > binom_table[16][26];
assign bits[16][27] = num > binom_table[16][27];
assign bits[16][28] = num > binom_table[16][28];
assign bits[16][29] = num > binom_table[16][29];
assign bits[16][30] = num > binom_table[16][30];
assign bits[16][31] = num > binom_table[16][31];
assign bits[16][32] = num > binom_table[16][32];

assign bits[17][1] = num > binom_table[17][1];
assign bits[17][2] = num > binom_table[17][2];
assign bits[17][3] = num > binom_table[17][3];
assign bits[17][4] = num > binom_table[17][4];
assign bits[17][5] = num > binom_table[17][5];
assign bits[17][6] = num > binom_table[17][6];
assign bits[17][7] = num > binom_table[17][7];
assign bits[17][8] = num > binom_table[17][8];
assign bits[17][9] = num > binom_table[17][9];
assign bits[17][10] = num > binom_table[17][10];
assign bits[17][11] = num > binom_table[17][11];
assign bits[17][12] = num > binom_table[17][12];
assign bits[17][13] = num > binom_table[17][13];
assign bits[17][14] = num > binom_table[17][14];
assign bits[17][15] = num > binom_table[17][15];
assign bits[17][16] = num > binom_table[17][16];
assign bits[17][17] = num > binom_table[17][17];
assign bits[17][18] = num > binom_table[17][18];
assign bits[17][19] = num > binom_table[17][19];
assign bits[17][20] = num > binom_table[17][20];
assign bits[17][21] = num > binom_table[17][21];
assign bits[17][22] = num > binom_table[17][22];
assign bits[17][23] = num > binom_table[17][23];
assign bits[17][24] = num > binom_table[17][24];
assign bits[17][25] = num > binom_table[17][25];
assign bits[17][26] = num > binom_table[17][26];
assign bits[17][27] = num > binom_table[17][27];
assign bits[17][28] = num > binom_table[17][28];
assign bits[17][29] = num > binom_table[17][29];
assign bits[17][30] = num > binom_table[17][30];
assign bits[17][31] = num > binom_table[17][31];
assign bits[17][32] = num > binom_table[17][32];

assign bits[18][1] = num > binom_table[18][1];
assign bits[18][2] = num > binom_table[18][2];
assign bits[18][3] = num > binom_table[18][3];
assign bits[18][4] = num > binom_table[18][4];
assign bits[18][5] = num > binom_table[18][5];
assign bits[18][6] = num > binom_table[18][6];
assign bits[18][7] = num > binom_table[18][7];
assign bits[18][8] = num > binom_table[18][8];
assign bits[18][9] = num > binom_table[18][9];
assign bits[18][10] = num > binom_table[18][10];
assign bits[18][11] = num > binom_table[18][11];
assign bits[18][12] = num > binom_table[18][12];
assign bits[18][13] = num > binom_table[18][13];
assign bits[18][14] = num > binom_table[18][14];
assign bits[18][15] = num > binom_table[18][15];
assign bits[18][16] = num > binom_table[18][16];
assign bits[18][17] = num > binom_table[18][17];
assign bits[18][18] = num > binom_table[18][18];
assign bits[18][19] = num > binom_table[18][19];
assign bits[18][20] = num > binom_table[18][20];
assign bits[18][21] = num > binom_table[18][21];
assign bits[18][22] = num > binom_table[18][22];
assign bits[18][23] = num > binom_table[18][23];
assign bits[18][24] = num > binom_table[18][24];
assign bits[18][25] = num > binom_table[18][25];
assign bits[18][26] = num > binom_table[18][26];
assign bits[18][27] = num > binom_table[18][27];
assign bits[18][28] = num > binom_table[18][28];
assign bits[18][29] = num > binom_table[18][29];
assign bits[18][30] = num > binom_table[18][30];
assign bits[18][31] = num > binom_table[18][31];
assign bits[18][32] = num > binom_table[18][32];

assign bits[19][1] = num > binom_table[19][1];
assign bits[19][2] = num > binom_table[19][2];
assign bits[19][3] = num > binom_table[19][3];
assign bits[19][4] = num > binom_table[19][4];
assign bits[19][5] = num > binom_table[19][5];
assign bits[19][6] = num > binom_table[19][6];
assign bits[19][7] = num > binom_table[19][7];
assign bits[19][8] = num > binom_table[19][8];
assign bits[19][9] = num > binom_table[19][9];
assign bits[19][10] = num > binom_table[19][10];
assign bits[19][11] = num > binom_table[19][11];
assign bits[19][12] = num > binom_table[19][12];
assign bits[19][13] = num > binom_table[19][13];
assign bits[19][14] = num > binom_table[19][14];
assign bits[19][15] = num > binom_table[19][15];
assign bits[19][16] = num > binom_table[19][16];
assign bits[19][17] = num > binom_table[19][17];
assign bits[19][18] = num > binom_table[19][18];
assign bits[19][19] = num > binom_table[19][19];
assign bits[19][20] = num > binom_table[19][20];
assign bits[19][21] = num > binom_table[19][21];
assign bits[19][22] = num > binom_table[19][22];
assign bits[19][23] = num > binom_table[19][23];
assign bits[19][24] = num > binom_table[19][24];
assign bits[19][25] = num > binom_table[19][25];
assign bits[19][26] = num > binom_table[19][26];
assign bits[19][27] = num > binom_table[19][27];
assign bits[19][28] = num > binom_table[19][28];
assign bits[19][29] = num > binom_table[19][29];
assign bits[19][30] = num > binom_table[19][30];
assign bits[19][31] = num > binom_table[19][31];
assign bits[19][32] = num > binom_table[19][32];

assign bits[20][1] = num > binom_table[20][1];
assign bits[20][2] = num > binom_table[20][2];
assign bits[20][3] = num > binom_table[20][3];
assign bits[20][4] = num > binom_table[20][4];
assign bits[20][5] = num > binom_table[20][5];
assign bits[20][6] = num > binom_table[20][6];
assign bits[20][7] = num > binom_table[20][7];
assign bits[20][8] = num > binom_table[20][8];
assign bits[20][9] = num > binom_table[20][9];
assign bits[20][10] = num > binom_table[20][10];
assign bits[20][11] = num > binom_table[20][11];
assign bits[20][12] = num > binom_table[20][12];
assign bits[20][13] = num > binom_table[20][13];
assign bits[20][14] = num > binom_table[20][14];
assign bits[20][15] = num > binom_table[20][15];
assign bits[20][16] = num > binom_table[20][16];
assign bits[20][17] = num > binom_table[20][17];
assign bits[20][18] = num > binom_table[20][18];
assign bits[20][19] = num > binom_table[20][19];
assign bits[20][20] = num > binom_table[20][20];
assign bits[20][21] = num > binom_table[20][21];
assign bits[20][22] = num > binom_table[20][22];
assign bits[20][23] = num > binom_table[20][23];
assign bits[20][24] = num > binom_table[20][24];
assign bits[20][25] = num > binom_table[20][25];
assign bits[20][26] = num > binom_table[20][26];
assign bits[20][27] = num > binom_table[20][27];
assign bits[20][28] = num > binom_table[20][28];
assign bits[20][29] = num > binom_table[20][29];
assign bits[20][30] = num > binom_table[20][30];
assign bits[20][31] = num > binom_table[20][31];
assign bits[20][32] = num > binom_table[20][32];

assign bits[21][1] = num > binom_table[21][1];
assign bits[21][2] = num > binom_table[21][2];
assign bits[21][3] = num > binom_table[21][3];
assign bits[21][4] = num > binom_table[21][4];
assign bits[21][5] = num > binom_table[21][5];
assign bits[21][6] = num > binom_table[21][6];
assign bits[21][7] = num > binom_table[21][7];
assign bits[21][8] = num > binom_table[21][8];
assign bits[21][9] = num > binom_table[21][9];
assign bits[21][10] = num > binom_table[21][10];
assign bits[21][11] = num > binom_table[21][11];
assign bits[21][12] = num > binom_table[21][12];
assign bits[21][13] = num > binom_table[21][13];
assign bits[21][14] = num > binom_table[21][14];
assign bits[21][15] = num > binom_table[21][15];
assign bits[21][16] = num > binom_table[21][16];
assign bits[21][17] = num > binom_table[21][17];
assign bits[21][18] = num > binom_table[21][18];
assign bits[21][19] = num > binom_table[21][19];
assign bits[21][20] = num > binom_table[21][20];
assign bits[21][21] = num > binom_table[21][21];
assign bits[21][22] = num > binom_table[21][22];
assign bits[21][23] = num > binom_table[21][23];
assign bits[21][24] = num > binom_table[21][24];
assign bits[21][25] = num > binom_table[21][25];
assign bits[21][26] = num > binom_table[21][26];
assign bits[21][27] = num > binom_table[21][27];
assign bits[21][28] = num > binom_table[21][28];
assign bits[21][29] = num > binom_table[21][29];
assign bits[21][30] = num > binom_table[21][30];
assign bits[21][31] = num > binom_table[21][31];
assign bits[21][32] = num > binom_table[21][32];

assign bits[22][1] = num > binom_table[22][1];
assign bits[22][2] = num > binom_table[22][2];
assign bits[22][3] = num > binom_table[22][3];
assign bits[22][4] = num > binom_table[22][4];
assign bits[22][5] = num > binom_table[22][5];
assign bits[22][6] = num > binom_table[22][6];
assign bits[22][7] = num > binom_table[22][7];
assign bits[22][8] = num > binom_table[22][8];
assign bits[22][9] = num > binom_table[22][9];
assign bits[22][10] = num > binom_table[22][10];
assign bits[22][11] = num > binom_table[22][11];
assign bits[22][12] = num > binom_table[22][12];
assign bits[22][13] = num > binom_table[22][13];
assign bits[22][14] = num > binom_table[22][14];
assign bits[22][15] = num > binom_table[22][15];
assign bits[22][16] = num > binom_table[22][16];
assign bits[22][17] = num > binom_table[22][17];
assign bits[22][18] = num > binom_table[22][18];
assign bits[22][19] = num > binom_table[22][19];
assign bits[22][20] = num > binom_table[22][20];
assign bits[22][21] = num > binom_table[22][21];
assign bits[22][22] = num > binom_table[22][22];
assign bits[22][23] = num > binom_table[22][23];
assign bits[22][24] = num > binom_table[22][24];
assign bits[22][25] = num > binom_table[22][25];
assign bits[22][26] = num > binom_table[22][26];
assign bits[22][27] = num > binom_table[22][27];
assign bits[22][28] = num > binom_table[22][28];
assign bits[22][29] = num > binom_table[22][29];
assign bits[22][30] = num > binom_table[22][30];
assign bits[22][31] = num > binom_table[22][31];
assign bits[22][32] = num > binom_table[22][32];

assign bits[23][1] = num > binom_table[23][1];
assign bits[23][2] = num > binom_table[23][2];
assign bits[23][3] = num > binom_table[23][3];
assign bits[23][4] = num > binom_table[23][4];
assign bits[23][5] = num > binom_table[23][5];
assign bits[23][6] = num > binom_table[23][6];
assign bits[23][7] = num > binom_table[23][7];
assign bits[23][8] = num > binom_table[23][8];
assign bits[23][9] = num > binom_table[23][9];
assign bits[23][10] = num > binom_table[23][10];
assign bits[23][11] = num > binom_table[23][11];
assign bits[23][12] = num > binom_table[23][12];
assign bits[23][13] = num > binom_table[23][13];
assign bits[23][14] = num > binom_table[23][14];
assign bits[23][15] = num > binom_table[23][15];
assign bits[23][16] = num > binom_table[23][16];
assign bits[23][17] = num > binom_table[23][17];
assign bits[23][18] = num > binom_table[23][18];
assign bits[23][19] = num > binom_table[23][19];
assign bits[23][20] = num > binom_table[23][20];
assign bits[23][21] = num > binom_table[23][21];
assign bits[23][22] = num > binom_table[23][22];
assign bits[23][23] = num > binom_table[23][23];
assign bits[23][24] = num > binom_table[23][24];
assign bits[23][25] = num > binom_table[23][25];
assign bits[23][26] = num > binom_table[23][26];
assign bits[23][27] = num > binom_table[23][27];
assign bits[23][28] = num > binom_table[23][28];
assign bits[23][29] = num > binom_table[23][29];
assign bits[23][30] = num > binom_table[23][30];
assign bits[23][31] = num > binom_table[23][31];
assign bits[23][32] = num > binom_table[23][32];

assign bits[24][1] = num > binom_table[24][1];
assign bits[24][2] = num > binom_table[24][2];
assign bits[24][3] = num > binom_table[24][3];
assign bits[24][4] = num > binom_table[24][4];
assign bits[24][5] = num > binom_table[24][5];
assign bits[24][6] = num > binom_table[24][6];
assign bits[24][7] = num > binom_table[24][7];
assign bits[24][8] = num > binom_table[24][8];
assign bits[24][9] = num > binom_table[24][9];
assign bits[24][10] = num > binom_table[24][10];
assign bits[24][11] = num > binom_table[24][11];
assign bits[24][12] = num > binom_table[24][12];
assign bits[24][13] = num > binom_table[24][13];
assign bits[24][14] = num > binom_table[24][14];
assign bits[24][15] = num > binom_table[24][15];
assign bits[24][16] = num > binom_table[24][16];
assign bits[24][17] = num > binom_table[24][17];
assign bits[24][18] = num > binom_table[24][18];
assign bits[24][19] = num > binom_table[24][19];
assign bits[24][20] = num > binom_table[24][20];
assign bits[24][21] = num > binom_table[24][21];
assign bits[24][22] = num > binom_table[24][22];
assign bits[24][23] = num > binom_table[24][23];
assign bits[24][24] = num > binom_table[24][24];
assign bits[24][25] = num > binom_table[24][25];
assign bits[24][26] = num > binom_table[24][26];
assign bits[24][27] = num > binom_table[24][27];
assign bits[24][28] = num > binom_table[24][28];
assign bits[24][29] = num > binom_table[24][29];
assign bits[24][30] = num > binom_table[24][30];
assign bits[24][31] = num > binom_table[24][31];
assign bits[24][32] = num > binom_table[24][32];

assign bits[25][1] = num > binom_table[25][1];
assign bits[25][2] = num > binom_table[25][2];
assign bits[25][3] = num > binom_table[25][3];
assign bits[25][4] = num > binom_table[25][4];
assign bits[25][5] = num > binom_table[25][5];
assign bits[25][6] = num > binom_table[25][6];
assign bits[25][7] = num > binom_table[25][7];
assign bits[25][8] = num > binom_table[25][8];
assign bits[25][9] = num > binom_table[25][9];
assign bits[25][10] = num > binom_table[25][10];
assign bits[25][11] = num > binom_table[25][11];
assign bits[25][12] = num > binom_table[25][12];
assign bits[25][13] = num > binom_table[25][13];
assign bits[25][14] = num > binom_table[25][14];
assign bits[25][15] = num > binom_table[25][15];
assign bits[25][16] = num > binom_table[25][16];
assign bits[25][17] = num > binom_table[25][17];
assign bits[25][18] = num > binom_table[25][18];
assign bits[25][19] = num > binom_table[25][19];
assign bits[25][20] = num > binom_table[25][20];
assign bits[25][21] = num > binom_table[25][21];
assign bits[25][22] = num > binom_table[25][22];
assign bits[25][23] = num > binom_table[25][23];
assign bits[25][24] = num > binom_table[25][24];
assign bits[25][25] = num > binom_table[25][25];
assign bits[25][26] = num > binom_table[25][26];
assign bits[25][27] = num > binom_table[25][27];
assign bits[25][28] = num > binom_table[25][28];
assign bits[25][29] = num > binom_table[25][29];
assign bits[25][30] = num > binom_table[25][30];
assign bits[25][31] = num > binom_table[25][31];
assign bits[25][32] = num > binom_table[25][32];

assign bits[26][1] = num > binom_table[26][1];
assign bits[26][2] = num > binom_table[26][2];
assign bits[26][3] = num > binom_table[26][3];
assign bits[26][4] = num > binom_table[26][4];
assign bits[26][5] = num > binom_table[26][5];
assign bits[26][6] = num > binom_table[26][6];
assign bits[26][7] = num > binom_table[26][7];
assign bits[26][8] = num > binom_table[26][8];
assign bits[26][9] = num > binom_table[26][9];
assign bits[26][10] = num > binom_table[26][10];
assign bits[26][11] = num > binom_table[26][11];
assign bits[26][12] = num > binom_table[26][12];
assign bits[26][13] = num > binom_table[26][13];
assign bits[26][14] = num > binom_table[26][14];
assign bits[26][15] = num > binom_table[26][15];
assign bits[26][16] = num > binom_table[26][16];
assign bits[26][17] = num > binom_table[26][17];
assign bits[26][18] = num > binom_table[26][18];
assign bits[26][19] = num > binom_table[26][19];
assign bits[26][20] = num > binom_table[26][20];
assign bits[26][21] = num > binom_table[26][21];
assign bits[26][22] = num > binom_table[26][22];
assign bits[26][23] = num > binom_table[26][23];
assign bits[26][24] = num > binom_table[26][24];
assign bits[26][25] = num > binom_table[26][25];
assign bits[26][26] = num > binom_table[26][26];
assign bits[26][27] = num > binom_table[26][27];
assign bits[26][28] = num > binom_table[26][28];
assign bits[26][29] = num > binom_table[26][29];
assign bits[26][30] = num > binom_table[26][30];
assign bits[26][31] = num > binom_table[26][31];
assign bits[26][32] = num > binom_table[26][32];

assign bits[27][1] = num > binom_table[27][1];
assign bits[27][2] = num > binom_table[27][2];
assign bits[27][3] = num > binom_table[27][3];
assign bits[27][4] = num > binom_table[27][4];
assign bits[27][5] = num > binom_table[27][5];
assign bits[27][6] = num > binom_table[27][6];
assign bits[27][7] = num > binom_table[27][7];
assign bits[27][8] = num > binom_table[27][8];
assign bits[27][9] = num > binom_table[27][9];
assign bits[27][10] = num > binom_table[27][10];
assign bits[27][11] = num > binom_table[27][11];
assign bits[27][12] = num > binom_table[27][12];
assign bits[27][13] = num > binom_table[27][13];
assign bits[27][14] = num > binom_table[27][14];
assign bits[27][15] = num > binom_table[27][15];
assign bits[27][16] = num > binom_table[27][16];
assign bits[27][17] = num > binom_table[27][17];
assign bits[27][18] = num > binom_table[27][18];
assign bits[27][19] = num > binom_table[27][19];
assign bits[27][20] = num > binom_table[27][20];
assign bits[27][21] = num > binom_table[27][21];
assign bits[27][22] = num > binom_table[27][22];
assign bits[27][23] = num > binom_table[27][23];
assign bits[27][24] = num > binom_table[27][24];
assign bits[27][25] = num > binom_table[27][25];
assign bits[27][26] = num > binom_table[27][26];
assign bits[27][27] = num > binom_table[27][27];
assign bits[27][28] = num > binom_table[27][28];
assign bits[27][29] = num > binom_table[27][29];
assign bits[27][30] = num > binom_table[27][30];
assign bits[27][31] = num > binom_table[27][31];
assign bits[27][32] = num > binom_table[27][32];

assign bits[28][1] = num > binom_table[28][1];
assign bits[28][2] = num > binom_table[28][2];
assign bits[28][3] = num > binom_table[28][3];
assign bits[28][4] = num > binom_table[28][4];
assign bits[28][5] = num > binom_table[28][5];
assign bits[28][6] = num > binom_table[28][6];
assign bits[28][7] = num > binom_table[28][7];
assign bits[28][8] = num > binom_table[28][8];
assign bits[28][9] = num > binom_table[28][9];
assign bits[28][10] = num > binom_table[28][10];
assign bits[28][11] = num > binom_table[28][11];
assign bits[28][12] = num > binom_table[28][12];
assign bits[28][13] = num > binom_table[28][13];
assign bits[28][14] = num > binom_table[28][14];
assign bits[28][15] = num > binom_table[28][15];
assign bits[28][16] = num > binom_table[28][16];
assign bits[28][17] = num > binom_table[28][17];
assign bits[28][18] = num > binom_table[28][18];
assign bits[28][19] = num > binom_table[28][19];
assign bits[28][20] = num > binom_table[28][20];
assign bits[28][21] = num > binom_table[28][21];
assign bits[28][22] = num > binom_table[28][22];
assign bits[28][23] = num > binom_table[28][23];
assign bits[28][24] = num > binom_table[28][24];
assign bits[28][25] = num > binom_table[28][25];
assign bits[28][26] = num > binom_table[28][26];
assign bits[28][27] = num > binom_table[28][27];
assign bits[28][28] = num > binom_table[28][28];
assign bits[28][29] = num > binom_table[28][29];
assign bits[28][30] = num > binom_table[28][30];
assign bits[28][31] = num > binom_table[28][31];
assign bits[28][32] = num > binom_table[28][32];

assign bits[29][1] = num > binom_table[29][1];
assign bits[29][2] = num > binom_table[29][2];
assign bits[29][3] = num > binom_table[29][3];
assign bits[29][4] = num > binom_table[29][4];
assign bits[29][5] = num > binom_table[29][5];
assign bits[29][6] = num > binom_table[29][6];
assign bits[29][7] = num > binom_table[29][7];
assign bits[29][8] = num > binom_table[29][8];
assign bits[29][9] = num > binom_table[29][9];
assign bits[29][10] = num > binom_table[29][10];
assign bits[29][11] = num > binom_table[29][11];
assign bits[29][12] = num > binom_table[29][12];
assign bits[29][13] = num > binom_table[29][13];
assign bits[29][14] = num > binom_table[29][14];
assign bits[29][15] = num > binom_table[29][15];
assign bits[29][16] = num > binom_table[29][16];
assign bits[29][17] = num > binom_table[29][17];
assign bits[29][18] = num > binom_table[29][18];
assign bits[29][19] = num > binom_table[29][19];
assign bits[29][20] = num > binom_table[29][20];
assign bits[29][21] = num > binom_table[29][21];
assign bits[29][22] = num > binom_table[29][22];
assign bits[29][23] = num > binom_table[29][23];
assign bits[29][24] = num > binom_table[29][24];
assign bits[29][25] = num > binom_table[29][25];
assign bits[29][26] = num > binom_table[29][26];
assign bits[29][27] = num > binom_table[29][27];
assign bits[29][28] = num > binom_table[29][28];
assign bits[29][29] = num > binom_table[29][29];
assign bits[29][30] = num > binom_table[29][30];
assign bits[29][31] = num > binom_table[29][31];
assign bits[29][32] = num > binom_table[29][32];

assign bits[30][1] = num > binom_table[30][1];
assign bits[30][2] = num > binom_table[30][2];
assign bits[30][3] = num > binom_table[30][3];
assign bits[30][4] = num > binom_table[30][4];
assign bits[30][5] = num > binom_table[30][5];
assign bits[30][6] = num > binom_table[30][6];
assign bits[30][7] = num > binom_table[30][7];
assign bits[30][8] = num > binom_table[30][8];
assign bits[30][9] = num > binom_table[30][9];
assign bits[30][10] = num > binom_table[30][10];
assign bits[30][11] = num > binom_table[30][11];
assign bits[30][12] = num > binom_table[30][12];
assign bits[30][13] = num > binom_table[30][13];
assign bits[30][14] = num > binom_table[30][14];
assign bits[30][15] = num > binom_table[30][15];
assign bits[30][16] = num > binom_table[30][16];
assign bits[30][17] = num > binom_table[30][17];
assign bits[30][18] = num > binom_table[30][18];
assign bits[30][19] = num > binom_table[30][19];
assign bits[30][20] = num > binom_table[30][20];
assign bits[30][21] = num > binom_table[30][21];
assign bits[30][22] = num > binom_table[30][22];
assign bits[30][23] = num > binom_table[30][23];
assign bits[30][24] = num > binom_table[30][24];
assign bits[30][25] = num > binom_table[30][25];
assign bits[30][26] = num > binom_table[30][26];
assign bits[30][27] = num > binom_table[30][27];
assign bits[30][28] = num > binom_table[30][28];
assign bits[30][29] = num > binom_table[30][29];
assign bits[30][30] = num > binom_table[30][30];
assign bits[30][31] = num > binom_table[30][31];
assign bits[30][32] = num > binom_table[30][32];

assign bits[31][1] = num > binom_table[31][1];
assign bits[31][2] = num > binom_table[31][2];
assign bits[31][3] = num > binom_table[31][3];
assign bits[31][4] = num > binom_table[31][4];
assign bits[31][5] = num > binom_table[31][5];
assign bits[31][6] = num > binom_table[31][6];
assign bits[31][7] = num > binom_table[31][7];
assign bits[31][8] = num > binom_table[31][8];
assign bits[31][9] = num > binom_table[31][9];
assign bits[31][10] = num > binom_table[31][10];
assign bits[31][11] = num > binom_table[31][11];
assign bits[31][12] = num > binom_table[31][12];
assign bits[31][13] = num > binom_table[31][13];
assign bits[31][14] = num > binom_table[31][14];
assign bits[31][15] = num > binom_table[31][15];
assign bits[31][16] = num > binom_table[31][16];
assign bits[31][17] = num > binom_table[31][17];
assign bits[31][18] = num > binom_table[31][18];
assign bits[31][19] = num > binom_table[31][19];
assign bits[31][20] = num > binom_table[31][20];
assign bits[31][21] = num > binom_table[31][21];
assign bits[31][22] = num > binom_table[31][22];
assign bits[31][23] = num > binom_table[31][23];
assign bits[31][24] = num > binom_table[31][24];
assign bits[31][25] = num > binom_table[31][25];
assign bits[31][26] = num > binom_table[31][26];
assign bits[31][27] = num > binom_table[31][27];
assign bits[31][28] = num > binom_table[31][28];
assign bits[31][29] = num > binom_table[31][29];
assign bits[31][30] = num > binom_table[31][30];
assign bits[31][31] = num > binom_table[31][31];
assign bits[31][32] = num > binom_table[31][32];

assign bits[32][1] = num > binom_table[32][1];
assign bits[32][2] = num > binom_table[32][2];
assign bits[32][3] = num > binom_table[32][3];
assign bits[32][4] = num > binom_table[32][4];
assign bits[32][5] = num > binom_table[32][5];
assign bits[32][6] = num > binom_table[32][6];
assign bits[32][7] = num > binom_table[32][7];
assign bits[32][8] = num > binom_table[32][8];
assign bits[32][9] = num > binom_table[32][9];
assign bits[32][10] = num > binom_table[32][10];
assign bits[32][11] = num > binom_table[32][11];
assign bits[32][12] = num > binom_table[32][12];
assign bits[32][13] = num > binom_table[32][13];
assign bits[32][14] = num > binom_table[32][14];
assign bits[32][15] = num > binom_table[32][15];
assign bits[32][16] = num > binom_table[32][16];
assign bits[32][17] = num > binom_table[32][17];
assign bits[32][18] = num > binom_table[32][18];
assign bits[32][19] = num > binom_table[32][19];
assign bits[32][20] = num > binom_table[32][20];
assign bits[32][21] = num > binom_table[32][21];
assign bits[32][22] = num > binom_table[32][22];
assign bits[32][23] = num > binom_table[32][23];
assign bits[32][24] = num > binom_table[32][24];
assign bits[32][25] = num > binom_table[32][25];
assign bits[32][26] = num > binom_table[32][26];
assign bits[32][27] = num > binom_table[32][27];
assign bits[32][28] = num > binom_table[32][28];
assign bits[32][29] = num > binom_table[32][29];
assign bits[32][30] = num > binom_table[32][30];
assign bits[32][31] = num > binom_table[32][31];
assign bits[32][32] = num > binom_table[32][32];

assign xorbits[2] = colbits[1]^colbits[2];
assign xorbits[3] = colbits[2]^colbits[3];
assign xorbits[4] = colbits[3]^colbits[4];
assign xorbits[5] = colbits[4]^colbits[5];
assign xorbits[6] = colbits[5]^colbits[6];
assign xorbits[7] = colbits[6]^colbits[7];
assign xorbits[8] = colbits[7]^colbits[8];
assign xorbits[9] = colbits[8]^colbits[9];
assign xorbits[10] = colbits[9]^colbits[10];
assign xorbits[11] = colbits[10]^colbits[11];
assign xorbits[12] = colbits[11]^colbits[12];
assign xorbits[13] = colbits[12]^colbits[13];
assign xorbits[14] = colbits[13]^colbits[14];
assign xorbits[15] = colbits[14]^colbits[15];
assign xorbits[16] = colbits[15]^colbits[16];
assign xorbits[17] = colbits[16]^colbits[17];
assign xorbits[18] = colbits[17]^colbits[18];
assign xorbits[19] = colbits[18]^colbits[19];
assign xorbits[20] = colbits[19]^colbits[20];
assign xorbits[21] = colbits[20]^colbits[21];
assign xorbits[22] = colbits[21]^colbits[22];
assign xorbits[23] = colbits[22]^colbits[23];
assign xorbits[24] = colbits[23]^colbits[24];
assign xorbits[25] = colbits[24]^colbits[25];
assign xorbits[26] = colbits[25]^colbits[26];
assign xorbits[27] = colbits[26]^colbits[27];
assign xorbits[28] = colbits[27]^colbits[28];
assign xorbits[29] = colbits[28]^colbits[29];
assign xorbits[30] = colbits[29]^colbits[30];
assign xorbits[31] = colbits[30]^colbits[31];
assign xorbits[32] = colbits[31]^colbits[32];

endmodule